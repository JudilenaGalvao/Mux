library verilog;
use verilog.vl_types.all;
entity MUX_vlg_vec_tst is
end MUX_vlg_vec_tst;
